`timescale 1ns/10ps
`include "define.h"
module test();
   reg[`BUS_ADDR_WIDTH-1:0] addr0;
   reg [`DATA_WIDTH-1:0]    idata0;
   wire [`DATA_WIDTH-1:0]   odata0;
   reg 			    rw0_;
   reg 			    breq0_;
   wire 		    bgrt0_;
   reg [`BUS_ADDR_WIDTH-1:0] dsaddr;
   reg [`BUS_ADDR_WIDTH-1:0] ddaddr;
   reg [1:0] 		     dmode;
   reg 			     dreq_;
   wire		     eop_;
   reg 			    reset_, clk;
   top u0(addr0, idata0, odata0, rw0_, breq0_, bgrt0_, dsaddr, ddaddr, dmode, dreq_, eop_, reset_, clk);
   always begin
      clk <= 1;
      #1;
      clk <= 0;
      #1;
   end
   initial begin
      #1;
      $dumpfile("dump.vcd");
      $dumpvars(0, test.u0);
      reset_ <= `Enable_;
      #5;
      reset_ <= `Enable_;
      #5;
      reset_ <= `Disable_;
      #5;
      
      addr0 <= 10'h150;
      idata0 <= 8'h99;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h150;
      idata0 <= 0;
      #2;
      $display("processor read and write");
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Disable_;
      dsaddr <= 10'h150;
      ddaddr <= 10'h160;
      dmode <= `Single;
      dreq_ <= `Enable_;
      #1;
      dreq_ <= `Disable_;
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h160;
      idata0 <= 0;
      #2;
      $display("DMA single mode");
      $display("addr = %h odata = %h", addr0, odata0);
      #5;
      addr0 <= 10'h151;
      idata0 <= 8'h98;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h151;
      idata0 <= 0;
      #2;
      $display(" ");
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      
      addr0 <= 10'h152;
      idata0 <= 8'h97;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h152;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      
      addr0 <= 10'h153;
      idata0 <= 8'h96;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h153;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      addr0 <= 10'h204;
      idata0 <= 8'h4;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      addr0 <= 10'h204;
      idata0 <= 8'h1;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      addr0 <= 10'h170;
      idata0 <= 8'h2;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h170;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      addr0 <= 10'h171;
      idata0 <= 8'h5;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h171;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      addr0 <= 10'h172;
      idata0 <= 8'h4;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h172;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      #2;
      addr0 <= 10'h173;
      idata0 <= 8'h2;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      
      #2;
      rw0_ <= `Read;
      addr0 <= 10'h173;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Disable_;
      dsaddr <= 10'h150;
      ddaddr <= 10'h160;
      dmode <= `BURST_MEM_MEM;
      dreq_ <= `Enable_;
      #1;
      dreq_ <= `Disable_;
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h160;
      idata0 <= 0;
      #2;
      $display("DMA burst memory to memory(from 150 to 160)");
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h161;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h162;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h163;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Disable_;
      dsaddr <= 10'h170;
      ddaddr <= 10'h204;
      dmode <= `BURST_MEM_IO;
      dreq_ <= `Enable_;
      #8;
      dreq_ <= `Disable_;
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h200;
      idata0 <= 0;
      #5;
      $display("DMA burst memory to IO(from 170 to 204)");
      $display("addr = %h odata = %h", addr0, odata0);
      #5;
      addr0 <= 10'h204;
      idata0 <= 2;
      rw0_ <= `Write;
      breq0_ <= `Enable_;
      dreq_ <= `Disable_;
      #5;
      breq0_ <= `Disable_;
      dsaddr <= 10'h200;
      ddaddr <= 10'h180;
      dmode <= `BURST_IO_MEM;
      dreq_ <= `Enable_;
      #10;
      dreq_ <= `Disable_;
      #5;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h180;
      idata0 <= 0;
      #10;
      $display("DMA burst IO to memory(from 200 to 180");
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h181;
      idata0 <= 0;
      #5;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h182;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #2;
      breq0_ <= `Enable_;
      rw0_ <= `Read;
      addr0 <= 10'h183;
      idata0 <= 0;
      #2;
      $display("addr = %h odata = %h", addr0, odata0);
      #5;
      $finish;
      
   end // initial begin
endmodule // test

   
